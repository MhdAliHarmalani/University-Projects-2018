PK     ! ߤ�lZ      [Content_Types].xml �(�                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                 ���n�0E�����Ub袪*�>�-R�{V��Ǽ��QU�
l"%3��3Vƃ�ښl	�w%�=���^i7+���-d&�0�A�6�l4��L60#�Ò�S
O����X� �*��V$z�3��3������%p)O�^����5}nH"d�s�Xg�L�`���|�ԟ�|�P�rۃs��?�PW��tt4Q+��"�wa���|T\y���,N���U�%���-D/��ܚ��X�ݞ�(���<E��)�� ;�N�L?�F�˼��܉��<Fk�	�h�y����ڜ���q�i��?�ޯl��i� 1��]�H�g��m�@����m�  �� PK     ! ���   N   _rels/.rels �(�                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                 ���j�0@���ѽQ���N/c���[IL��j���<��]�aG��ӓ�zs�Fu��]��U��	��^�[��x ����1x�p����f��#I)ʃ�Y���������*D��i")��c$���qU���~3��1��jH[{�=E����~
f?��3-���޲]�Tꓸ2�j)�,l0/%��b�
���z���ŉ�,	�	�/�|f\Z���?6�!Y�_�o�]A�  �� PK     ! �d�Q�   1   word/_rels/document.xml.rels �(�                                                                                                                                                                                                                                                                 ���j�0E�����}-;}PB�lJ!��� E?�,	��`HI��`��r��sπ6����w��{���r茯{�*x���AkWk�*�`[^^l��jNK���D�8R�1���d:4e>�K/����4�Vm^u�r��w2NP�0ŮVw�5�j��o����7o:>S!?p����8JX[d�0KD��EVK���c2�P,���ũ�a���]���.���ﰘs�Yҡ�+�����(!O>z�  �� PK     ! 
_���  �J     word/document.xml�\[o�8~_i����i�����aVӖ�"ͥ�e��d'XM��1P���q�@!$��� Ď��9߹96|����P���rV�̊�!�,nS�ֵۛ���3{���6$��O��>j6�z>a	��U׺R5]�.�qX�%x�Y���sǡ�\���aѷ@p��!�w�Y�ZBκOG�x ���nu���~B�\�ȑ�Q?�%�ϋ� ����.���X���2����Q9����k=�j	��5���|�F�4��C�8�uA<����K��N��Ԡ�;"�_$D��F����A�ǨL�a?���b�S4��(�iX��sĉ�)�L�I5�k�F�`��qHV#q���á?q�Aஇ��`B��G���ƴT�Z�Vb--8\���.��}��r��G�=�P� R^�5 �v�=T�� �Wu�0�?~��4��<9�s��)""8w�B@�0�+�-!�i���M6<�X?��B�G�n2��P��Z`�AB"�Dk�V���4Eރ���|E�\ߜ����h��M�Z�������U����/����ŏ�y��F<墯Dex�[(�����]��y\�5�84���a �:�2U�I
�-�E���N�`�c���2v�A}*i���P"��R�r@#�n��[�t��p�_-�#���s^�u�.,
�=��R����^��FA	P��g���m��|yN�'x��fl���1l�#K�$���P�{2G<�$��j����B��Yy���I�#sFiCMYK��f/ض�X�j����G�B;�VA�	]D;΄-
+h�(k)��'\/nZ�bF���+�/�6Bi�=�R+�`E�PK����)��������%Y�V��+����p={�z�լ����TK�D�sNI�)�C�y3+��*W}7,�����\�a�j�@�#��ְ�qΟ�mZ��-�!u^��(�iٗ��(��!5��P��,����s�'��ahOW��s1�o�Ii��a���8;0����Fu���p(�`�E�/�KN�w��o����l�(���E��s���fO�`+Ʃ�9�a]HSʅ;�]"�l��pO�Kh�-:ĥl�s�1b�I�x(�3n����e�7�i�0���>+�w;�����n���w�f#y��j+7#G�R1~]��lYtX�G���L�����=u uZ�\e��g�rX�c��\U��t�B����Γ�y)�Ju��V�s�#��oNo+�5��5�K���h�@���
�����#�n�.s=��21T.K�||GP����l���A��Ȧ�X�Ng�U�_S��.-RBJ�py�����E�ZՌʇ��K�+:U��62�PC�>ay���ގ��	��9��5
Aq�_'Q�,?g�6e��$�#ht���P��,:3���:/����=#�*sˣ`��	I�4���Xl�{���V��C�T��H,��T{�����t-�%����䠢��nٖM#c\����	���hٱ�+Y�����2��2�J=���wxA�܄e��b�~9><��2Ě�J������_E ej��u�}�Ѿ�غ���s�<�NH,y���UQļ{��u�<8�F3t���I5��n��#�x ���Aݮ�\v��ܟ\{�y�ۅe2u��At�p.\�=]&�Y��5Q��'j��u!�ϣ�\Ri���#9c���_���j�  �� PK     ! �@�$  �     word/theme/theme1.xml�YM�7����;�3�X�㱝��MBv���<#�(֌�$�	���z)��C��PJ4����Ц?���c�l�K���5������H�z�,��	���k׮8���D(�����a�m[��,�d�k�!�����U���BK�glt���^��B��2����.�4�F�
�)���YM�l+�p{{<F!���K{�p>��_ƙl1=���f��Ѥ&�؜�Z' wm1NDN���-]�Qvu�jui��ے�P�-�Ѥ��h<Z���6���|7h���ҟ�03͹��^���{l	����~���K�xߓ�@y�����*�%P^�1i�W�+P^ln�[��w[^�����񚍠��2&�����a����P�����3�m���!�CP�e�O�� �FY(N���0��ԝ�����U%�A�:o
�F��c���)�ڟ
�v	��ի�'/ϟ�z������co�� Y\�{��W=������>�ڌge����x�����k��y�����~�Ǐ�p��Q~�RȬ[�ԺKR1A� pD���8�l�g1�6�'��``�����Tȅ	x}�P#|��G��$Հ�����9ݔc��0�b��tV����4v����l*�=2��Ѽ�E�A3�-�G&� �����02��d� 2����մ2��R�����ȷ���V�`��><ёbo lr	���`�AjdR\F ��H�i��q��bb"Ș��6�kto
�1���SI9�����2�O&Aҩ�3ʒ2�6KXw7� ��u��mM�}�t_���	2/�3��-���x�r^]��e����{�Oޅ����Ysw �f�e�ܧȸ��%|n]�B#���v̲;Pl���_���m?�^�W��.��u]�I�����#>���)egbz�P4��2Z>*LQ\��b
T٢��xr�����F���u̬)a�lP�F߲��C孵Z�t* _����h'�[���c�ҽ���q�  m߅Di0�D�@�U4^@B�l',:m�~+��Ȋ��?lxn�H�7�a$����y��S�v�0��些Lk$J�M'QZ�	��z�s�Y�T�'C�I��~��"��8�k֩�sO�	��k�ŭPө�Ǥng];�@�e�R���%9Lu��O���(k�������-9��\���"���I��1���UU��N����
�	�GItj����"P^�&!Ɨь--�U��j��_�V[�i'JY�s�*/�桘��J�/&3�e�.}�^l$;J��� ���Y?��!_b��}�U.��Z�)�n�)q��Dm5�FM26P[���vx!(�\��Έ]��VŽR�6^O��C����:Ü)��L<#�˹��B]θ5��k?r<��^Pq�ޠ�6\����F���Fm�՜~��X�'i�����<_�}Q�o`��}%$i��{pU�70���70�yԬ;�N�Y�4�a���ڕN��U�͠����>��v�F�6�J���H��N������������y�]�W���  �� PK     ! ��&�  %
     word/settings.xml�V�n�8}_`�A��*�|�P���x�"�.*�(�������.��wH�����E�L͙93$����gўhC����UGD�S��ǟ7�dG�"�����#1���{{(��L����;kU�����̕TD �H͑�O�M9ҏ�Jj������c:ȲI���y�jQ�	���F6օ�ihM���/�ۅ,e�r"�Ϙj )̎*���epH���Ğ��wȳ�{�?G\R�PZ��� �B�T��^=羂��=��_�W>�1��+��!?F1�)Rs��)vɑt��4ҝ����uq�R��A9p.l-���נ�/R��P(�k�jh�,�S�˦����"����A@{(�qP{��L�2�AUi��=�꧃���!�jKt�Pl�RX-Y���/io�s4\l���*����8��E��%&��V�������<�׉$�M1ٸs,푑_�/�F���}��D�+���#���Ȋ ��1��d�&V��5�Z�{�A�,m�!��A>T˃?��a�?�7=�<؄�')mpͲ�b0N�Jz	����o���M�oV>&}��7D��a�$�.��JS�ݘM�G�T�"���)�*�I��#�V�c���L�Z�Ư��퉷��ߴB?x�r��?�lU�4R�4�K>��T�ʃݴU��3���^�s:ϡ�pž�����%"�\�˭(9 ��7���.�*�)Չ��������.�����T�A�<6�0��j�Q��'� �����6<�F�6:���6>�&�6q�����:Kgo$c�@�������!E�������d���`j�?����'7�^��7CG���s��%F�{��U-�i�)��<��4��50<V���|�_�Q?��~"��{������'��r�'�E�LF��(�-�$��,ǫ����n�oߔ����   �� PK     ! �1��  D     word/fontTable.xmlܓ]k�0���B��e磝�Sڬ���E�~��ȶ�>��7�~ǒ��B���`�AH��y|�Z����h�����'�i��*�T������n�vVV� �>,?~����� �-�FT��+�D+����`������?vݍp��Am�V��-���VB~vbg�1?�R#�YhUGZ�Z����NH <�щg��'L>;%�W�	f�(�0=gqf�/��:@qX��1�|�Ĉ�Kc���$<��H���3I_Zn0��Zm����[2�؞늲����᝱�0�l�(Z�A��q�Jr͍҇�
�H�N��=�j(-�@5���U��1V<��4)9�ev�4*��O�2=)lPD��e�8"rN{�Yr�̉G,K_��-Ё�Dt�������w��ë2�7ٓg���H��L�v���^刏�Ǒ�G�Wմ�b���v�8��O   �� PK     ! �?�b"  N     word/webSettings.xml���J1 ��;���l�-�t[����{�ζ�$2����תH/�-��|�$��vމwHd1Tr�/��`peú���y�R
�:��� �l��lz~6i��ϐ3�$�J�қJnr��Rd6�5�1B�d����aZ+���6����]Zgs��E1�{&�`][�h�B��U�"��H?Zs��`Zń�x�=�m�e��&!a��<̾����Aѭ��F��`Lp1��Z;)�)o��^:�x$�]��S~R��z�sLW	�����^���z�E�9l�n8P�~��  �� PK     ! ���x  �   docProps/app.xml �(�                                                                                                                                                                                                                                                                 �RMO�0�#���Y�M �� 4�8�%�l�(qۈ4��l��=�2'r�������7�C��.��*��)m�E�Zߝ]�EL�*a��Ey�X^��x	�cHcA6.�.%�X��"N�l�ҸЋDih�k-���m�6�YU]0�'�
ՙ	ˁ�j��K�����>x��Pc�Hȟ�(�z`#
�K�ԺG^<&�"Z�|
l`り|6�6���D2��|:���� ���h)���.�&���L �h��m�鐅��m�B��� � |�<3XIapI�F����X��K|l���-����f/>G~�Gknt�V^�,�<�g	V���F# ��*��hֶ��z~����{��Ť����F�����  �� PK     ! ���r  �   docProps/core.xml �(�                                                                                                                                                                                                                                                                 ��MO�0��H��*�6i���N|h��$$�@�B�mai%���=i�vT��͎�v�$�}�2؃��R9�#�P��B�s����7(��*Ne� G�hV\^dL��2�l*�	��WR6e:G�t��e(��<�|qU��:��5֔m�pB�5.�QNō`�Et��l��;#[�0H(A9��(�'ց)�ن��,�;h8��Ł��b 뺎�I���c��xzi�
�x� g�NB��S�#�����!�13@]e�ņ�J<RJ�`_ll�¡��^b�y��eFh��0:��-���ÙY����^4?���ĐfG����ަ�3���M��sT$$!!���tI��8N	�hV�����V�:��_��  �� PK     ! ��*  Sp     word/styles.xml��]sۺ��;����U{���g�9�ۉkO���i�!�P��ʏ��/ R�%(.���-Q� ċ������ϩ�~�*;M��"��*������ջ��(Y�0�2~6z����O��oO�E�"yi@V����hQ����<e�{��>8Wy�J�2�,���b�.Y)fB��e���w<j0y���E�?��JyV��qΥ&��X�e��=��=�<Y�*�E�O:�5/e"[c&� ��8W������45�(>ٳ��r8����8�Q�/)Ei|z󐩜ͤ&�S�t�"}�j&*��笒ea^�wy�ye�\��,��SV�B��ZhT*4��<+�H�(��Z.�?�G�t޾��M����_L����W�\�l�'Y��z�g�~Lݚ8o�4�l��w�s8nN������+[����%�ur�g�R_�}\��^�fU��B,���ƎA����{�6�>��_U�ȓi���lY��7w�P�6���-S�9婸I�3��B$��g?
�l����v��XU����db{�,�/�1_+�3�|3�|���m�V�I�D[��33�D��[}b�D�ٶ3�W�n?�*��
:|���ު��*��
��VY��� �%��6",Pwq<nDs<fCs<^Bs<VAs<N@s<���c4��M�Rž^�t�Oo���#¸���0�� ��{����ø���0���;��{��s�Vt�m���]6W��Tɣ�?��L�l�E�3��IN� S�l�D<�3�zw�&��K��Ej��C���|h�y��K�%G,I4����=-ҧs>�9�bNٱ�&��*���%{ c�,!n��dPXwh�?/�IA�NY���US�l|�*��me �E%%'b}��b�5<7��ᩁ��,fxb�hF�D���Q�54�v��'U�54�vkhD��І�۽(���UǤ��ݥTf[|p=��!cz0|�i�L�;����-�ٕnǺ�-�B%/�=Ŝ�&Q��m��g-�jx�nѨ̵��k�#2ؚ7�b�z�lh�4�̴������^��2Y���nc���1���2�c	z�7��5rR�|�Z�؆5�V�G%��5H�ZJ?���/K���q0�JI��xBG������k�}+I/�I�V�+m!�O����-[>�;�DF�ۗw)2�[A\��~���Ҥ��ah��,UJ�lv�����NS�s�g/Dg{N�=da��`��I*!"�e���jy��/3��v������,]֋o�q�I�?�!��˅��2�=	��6,�ٿy<|���"���?���?ڥ����_&l�/��zz0���d�p�OvGu�����^B�Q��G}�Ó�����畤k���W@�&T�J���-���-��|	���l�Y�?r���aaTJX�F����
0�6�66�^�F�p`T��t�'��������Q�3��gF��>G|>׋`�)�AR�9I7�d%O�*g����`�����jnnPY}7��QK��v���'��UͰ(�E�#ʤT�hom3����{�v��'9W�N��/�Lx�9'�Η��c��o��k��xX��t���w1�{;#W	�V�����x�<K[�-OD��*
�8>�l{�V�����Jb+�g$,�xw�f��y�3���g���Vd�>����#�t��u���|']�h�ZlWGZG�u���^�e��<����N?�������q��������W~D����_���AӖ��{��v�k���R������u��SV�s�����(�o��Í�{��#z@~D��������c��{��#У�p��ǍV0>d�����j�*����#�F��Q���QAx�Q!mT�@"�F�0�Qa<Ψ0>Ĩ�bTHA"�F��Q!mT�@5pm�2*���
h�Bڨv�8��0gTbTH	1*���
h�Bڨ�6*D��
(��� �B
ڨ�6*D��Z?jnT�3*�1*��R�F��Q!mT�@"�F��QAx�Q!mT�@"�F���
�C�
)!F��Q!mT�@"�F��Q!eTdTHA"�F�����\���f?��zz���骩�w�Qnu�������Y����l��"fR(�E��r�-��\v?���~�R�,��f
��}#���aW�w#A�w����H��<�}�H0v�֗��R�t���'x�	���p��]c�[�kdvaw��N�Qd���G=��x}) tuG�p�'tuK��j8���+���W=?���~JO//��V؏
��+u�Q��Ԑ$5��KQ�RCT��p`�J	X��g?!Hj�	������0��T���RCV��.5DKQaR��VjH�J	X�!!Hj�	������0�A����RCVjH�`¥��`�!�Kj���%5Ja'�sq������lɉ̖B`��Zi�˖\������	}e�Pzz1xa�(��~T�Ըl�M�p��	X�qْWj\��)5.[��-���eKmR㲥6��g?!Hj\��)5.[��-���eKmR㲥6�q�R��'d/&\j\��)5.[�K�˖ڤ�eKmR㲥6�qْWj\��)5.[��-���eKmR㲥6�q�R�Ըl�+5.[��-uJ�ɖ�O[?�d�����˗%7���<0���A�\��I�?�d�MM��'���m���u�6/tYq��I���oA]?�c��u���J��4���M�n.�֟ۺ��Y��4yG��$�mT���Ǧ��L�?ڥ���xj~���i��j�>~ɥ�e�����Q��e}t�g�u|V��7>��0ޮL����0O{���\��vI㆖涷Sm�M�V���  �� PK-      ! ߤ�lZ                      [Content_Types].xmlPK-      ! ���   N               �  _rels/.relsPK-      ! �d�Q�   1               �  word/_rels/document.xml.relsPK-      ! 
_���  �J               �  word/document.xmlPK-      ! �@�$  �               �  word/theme/theme1.xmlPK-      ! ��&�  %
               9  word/settings.xmlPK-      ! �1��  D               2  word/fontTable.xmlPK-      ! �?�b"  N               .  word/webSettings.xmlPK-      ! ���x  �               �  docProps/app.xmlPK-      ! ���r  �               0   docProps/core.xmlPK-      ! ��*  Sp               �"  word/styles.xmlPK      �  0.    