PK     ! ߤ�lZ      [Content_Types].xml �(�                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                 ���n�0E�����Ub袪*�>�-R�{V��Ǽ��QU�
l"%3��3Vƃ�ښl	�w%�=���^i7+���-d&�0�A�6�l4��L60#�Ò�S
O����X� �*��V$z�3��3������%p)O�^����5}nH"d�s�Xg�L�`���|�ԟ�|�P�rۃs��?�PW��tt4Q+��"�wa���|T\y���,N���U�%���-D/��ܚ��X�ݞ�(���<E��)�� ;�N�L?�F�˼��܉��<Fk�	�h�y����ڜ���q�i��?�ޯl��i� 1��]�H�g��m�@����m�  �� PK     ! ���   N   _rels/.rels �(�                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                 ���j�0@���ѽQ���N/c���[IL��j���<��]�aG��ӓ�zs�Fu��]��U��	��^�[��x ����1x�p����f��#I)ʃ�Y���������*D��i")��c$���qU���~3��1��jH[{�=E����~
f?��3-���޲]�Tꓸ2�j)�,l0/%��b�
���z���ŉ�,	�	�/�|f\Z���?6�!Y�_�o�]A�  �� PK     ! �d�Q�   1   word/_rels/document.xml.rels �(�                                                                                                                                                                                                                                                                 ���j�0E�����}-;}PB�lJ!��� E?�,	��`HI��`��r��sπ6����w��{���r茯{�*x���AkWk�*�`[^^l��jNK���D�8R�1���d:4e>�K/����4�Vm^u�r��w2NP�0ŮVw�5�j��o����7o:>S!?p����8JX[d�0KD��EVK���c2�P,���ũ�a���]���.���ﰘs�Yҡ�+�����(!O>z�  �� PK     ! �y�	  9     word/document.xml�[mS�8�~3�v�/7�ئ�rn��f�����J�C�<�����[��z�46C��ز��h���J&�>\�&Ti&E���Pɘ�q�1�l�6@"b¥��ƌ�Ƈ����n�2�S*���i��1Y�y:JhJt+e��Z�L+��'G#Qo*U�m���2%#�5�; bBt�]�OZ��;[��^�e��RF��Bv���ݛ����Ɍ
|8�*%o��K��̳&�͈aCƙ��H��\�l7r%�RDs�v	(�yu�E�N9N��(GR�e��?*&s!�ob���{�,�~�Ct�YY
��r*S^ �����ǌX���p]�IJ�X*�!Ӭ7��>[k^k�}"vJ����Иf���'%�l)�=LZW\.dY��Y���z�~��d�iv�B*2��p��� �(i�G6�xf�f0���v�G�o:�HeS��H����ӕ&+Dٓy����;�J�g���Ol��Dh�LQMՄ6pp`)U�B�4��P���T�(�b<�C��� ����Ý]@N��F�ݭm^;T����:hUX�X�9���7@<�K,q<tid��_g��#t�.4���3T��5I�*��*�/���5$��X��158q�7?ew�rQ��:���D�e�ت��Q�K���s}��UBRRK�t�� H]|�sw=w�zQDݓ�M�b%�Y�O����߆]	r���@>2d���п���6�
�K���n���t"1�USh����ԡ#��hR*��F�b�E�����ʱLnkj0��j�&��r�" �?X(��`RF��dg
�TF���\0���*7��?�3q�F�{b]X�c���0�S2��E#�%�ر�ir:��^ώ�@\�dL .e�����qN���xV�e�8�!1DR�u�
�)fD�&K3Nm��m�J�Y�4/v]l��U�ҟ{l�Qw�l��0J�ۍk`Mb5�����[{GG�VΉ6g�P4>%c�������W�Q�PL#ɹ��a��P5���8Ɯsa6*�
\D1��)F����%F�I��	�j ,1����VA��yJ:�Q�S������/�d,�+��)�=U�ޮv���s�x��bJNȄ��>._����Q��Ia����B�Je`��+�����`��˙�w|�;�0}D�k��w�Q�zw�3u!tO`�\�
b9X!�/�b���˛(�D�uoT��Y+���m�#�F�WL\�u��«�<6�.��F����*�7�]��f�� l�K�
�}+!l���Rih?����^����[n� Jĵ!X��5��wɰX��¡����7�������:�o:?VH%p�et	.$e��n_�>/�P�!Xoc�^��B0,�6H�~�+���Oݓ':�"�n1����c[F乹�C�[P���)Խ�X$�"��w֍�f�^Վf-��n6׎�f�)`�h�䦲p���7�Ǒ�l�+��Em`�t�D%I��~��j��񌛷����dJ0�-�e	�mՊh�6��h�;���x�O�*��ύ�D��%k�M�@#��CY������1��H�m6�'1�~@U�v�Ԫ�)ʢ��V�����u����
�]�Y�$?2�������2O-V�6xʙm=�l������p~3t�R^���#��b�j���/>�}]P�����os�ƫidN�-p�0��_�Ѵ�������wv����1���̰}�xE�qb��Ci�L����V�&� ��o���HJ�r;΍�-�E�kl-'־�c}R��3AO�����qCt��o�����  �� PK     ! �@�$  �     word/theme/theme1.xml�YM�7����;�3�X�㱝��MBv���<#�(֌�$�	���z)��C��PJ4����Ц?���c�l�K���5������H�z�,��	���k׮8���D(�����a�m[��,�d�k�!�����U���BK�glt���^��B��2����.�4�F�
�)���YM�l+�p{{<F!���K{�p>��_ƙl1=���f��Ѥ&�؜�Z' wm1NDN���-]�Qvu�jui��ے�P�-�Ѥ��h<Z���6���|7h���ҟ�03͹��^���{l	����~���K�xߓ�@y�����*�%P^�1i�W�+P^ln�[��w[^�����񚍠��2&�����a����P�����3�m���!�CP�e�O�� �FY(N���0��ԝ�����U%�A�:o
�F��c���)�ڟ
�v	��ի�'/ϟ�z������co�� Y\�{��W=������>�ڌge����x�����k��y�����~�Ǐ�p��Q~�RȬ[�ԺKR1A� pD���8�l�g1�6�'��``�����Tȅ	x}�P#|��G��$Հ�����9ݔc��0�b��tV����4v����l*�=2��Ѽ�E�A3�-�G&� �����02��d� 2����մ2��R�����ȷ���V�`��><ёbo lr	���`�AjdR\F ��H�i��q��bb"Ș��6�kto
�1���SI9�����2�O&Aҩ�3ʒ2�6KXw7� ��u��mM�}�t_���	2/�3��-���x�r^]��e����{�Oޅ����Ysw �f�e�ܧȸ��%|n]�B#���v̲;Pl���_���m?�^�W��.��u]�I�����#>���)egbz�P4��2Z>*LQ\��b
T٢��xr�����F���u̬)a�lP�F߲��C孵Z�t* _����h'�[���c�ҽ���q�  m߅Di0�D�@�U4^@B�l',:m�~+��Ȋ��?lxn�H�7�a$����y��S�v�0��些Lk$J�M'QZ�	��z�s�Y�T�'C�I��~��"��8�k֩�sO�	��k�ŭPө�Ǥng];�@�e�R���%9Lu��O���(k�������-9��\���"���I��1���UU��N����
�	�GItj����"P^�&!Ɨь--�U��j��_�V[�i'JY�s�*/�桘��J�/&3�e�.}�^l$;J��� ���Y?��!_b��}�U.��Z�)�n�)q��Dm5�FM26P[���vx!(�\��Έ]��VŽR�6^O��C����:Ü)��L<#�˹��B]θ5��k?r<��^Pq�ޠ�6\����F���Fm�՜~��X�'i�����<_�}Q�o`��}%$i��{pU�70���70�yԬ;�N�Y�4�a���ڕN��U�͠����>��v�F�6�J���H��N������������y�]�W���  �� PK     ! +��k�  �	     word/settings.xml�V�n�8}_`�A��*��	�:�c�����D�&@Rv����)1r��p[��Ԝ�q���o�>q��T�y�\�a@D-1�y�y����@$0bR�yx$:|{��o�&ƀ����9���Θ6�Lt�#��`#G>�vz�ڨ��E�V�Qs��q<7rvJ䃋��ZI-cMr�4�&Ï�P���M
Yw��"Na��zG[�����;��{μ�!�ϸ�A*�lqNz֠U�&ZC�8�	R1�^9z�}��+:W`���t�������4�1���D9y�4;�$=�@+�TO�����B*T1H����]x,�"%yKT����pbL�1�AUid*{�\�\�B�!�lQ]XJa�d^��Y�(h�`�fb<��|��@r{13k�a y���E�.z2=�u 	�@QL6�&�92���K��,~�iC����_��{	a#�.n�-Yd:(�o
�:�b�]S�����ۂѦ!
Pd��C�<�:�#��Ÿ�S�R��>Ii�j�Y\�e}�=I��z�-$�����!���v!~T�d)��b�x�(
�veN�F�o��xE`t�)Rv���4G��`�<���� �;�5R���)�y~����:Q+ٵ=zP���U�,,�0�{���[	X6'P'���ru�s��؍�rTq�DD�K�܊b�RQ���TiYA֨m{rU�d2�ݙĚ���к�j�X갴����EA{8����N�.��r�e^�����MG���fV���V��G�?Zy#��ߍ�+Q_�C-)�l��`��:���	�5������b����Nm���3/t-f�ۗ02�O�c���r�OCM���W�ƿ�gT�Vh�q0Ry�/�%S�j�����4�H<`X��ؾN�Ϳ�x��WwEt��Q�&Yt{Y�rZ,�b�,����a(����  �� PK     ! �1��  D     word/fontTable.xmlܓ]k�0���B��e磝�Sڬ���E�~��ȶ�>��7�~ǒ��B���`�AH��y|�Z����h�����'�i��*�T������n�vVV� �>,?~����� �-�FT��+�D+����`������?vݍp��Am�V��-���VB~vbg�1?�R#�YhUGZ�Z����NH <�щg��'L>;%�W�	f�(�0=gqf�/��:@qX��1�|�Ĉ�Kc���$<��H���3I_Zn0��Zm����[2�؞늲����᝱�0�l�(Z�A��q�Jr͍҇�
�H�N��=�j(-�@5���U��1V<��4)9�ev�4*��O�2=)lPD��e�8"rN{�Yr�̉G,K_��-Ё�Dt�������w��ë2�7ٓg���H��L�v���^刏�Ǒ�G�Wմ�b���v�8��O   �� PK     ! �?�b"  N     word/webSettings.xml���J1 ��;���l�-�t[����{�ζ�$2����תH/�-��|�$��vމwHd1Tr�/��`peú���y�R
�:��� �l��lz~6i��ϐ3�$�J�қJnr��Rd6�5�1B�d����aZ+���6����]Zgs��E1�{&�`][�h�B��U�"��H?Zs��`Zń�x�=�m�e��&!a��<̾����Aѭ��F��`Lp1��Z;)�)o��^:�x$�]��S~R��z�sLW	�����^���z�E�9l�n8P�~��  �� PK     ! *zC9~  �   docProps/app.xml �(�                                                                                                                                                                                                                                                                 �R�N�0�W���Yg�*Eh֨�� i��ٲ'�UǶl�ؿgLJ����4����ދ��}4����ݖ�UUh�S���򥽻�.���U�8��򌱼���98�!i�Qظ-���cQ8�����I��(��g��Ľ��#���j�'�
ե�	ˉ��-�/�r2���쉏C��7"!ʛf�\��(�.	��yE�����1�5����*�6��D2Q����k` ~xo����Z]������L ly���k�霅,[x�6K�l�H[}~�|���0�� x'LD` ع�K|l���W|���,~��.l�t^H�Po�fix1������a���J0�ڵ=��3�r���y�u������#���   �� PK     ! v�>r  �   docProps/core.xml �(�                                                                                                                                                                                                                                                                 ���O�0��M�Hߡ�1X�����8�񭶷�J�vC�{&qO���>���M��e�@Q��AHVq!7z]-��K%�E%!C4�//R�Vix֕m�)I�0����*�ذ-�������tI�K�+�vt8"��`)���V�W�":Jr6J��.:�0P���A�O�]��]�Y
�(8�ő�6b��C��!~_>�tW��l�b���
[@��S�"���f��1q1�@m�����{�έ�JсC��}M]in��$sôP�=f?`r���t����3��2m���hHwĘ�G����{Φ�7u������#���h�"WI'�|�+N�O��q�+�Kӯ��   �� PK     ! ��*  Sp     word/styles.xml��]sۺ��;����U{���g�9�ۉkO���i�!�P��ʏ��/ R�%(.���-Q� ċ������ϩ�~�*;M��"��*������ջ��(Y�0�2~6z����O��oO�E�"yi@V����hQ����<e�{��>8Wy�J�2�,���b�.Y)fB��e���w<j0y���E�?��JyV��qΥ&��X�e��=��=�<Y�*�E�O:�5/e"[c&� ��8W������45�(>ٳ��r8����8�Q�/)Ei|z󐩜ͤ&�S�t�"}�j&*��笒ea^�wy�ye�\��,��SV�B��ZhT*4��<+�H�(��Z.�?�G�t޾��M����_L����W�\�l�'Y��z�g�~Lݚ8o�4�l��w�s8nN������+[����%�ur�g�R_�}\��^�fU��B,���ƎA����{�6�>��_U�ȓi���lY��7w�P�6���-S�9婸I�3��B$��g?
�l����v��XU����db{�,�/�1_+�3�|3�|���m�V�I�D[��33�D��[}b�D�ٶ3�W�n?�*��
:|���ު��*��
��VY��� �%��6",Pwq<nDs<fCs<^Bs<VAs<N@s<���c4��M�Rž^�t�Oo���#¸���0�� ��{����ø���0���;��{��s�Vt�m���]6W��Tɣ�?��L�l�E�3��IN� S�l�D<�3�zw�&��K��Ej��C���|h�y��K�%G,I4����=-ҧs>�9�bNٱ�&��*���%{ c�,!n��dPXwh�?/�IA�NY���US�l|�*��me �E%%'b}��b�5<7��ᩁ��,fxb�hF�D���Q�54�v��'U�54�vkhD��І�۽(���UǤ��ݥTf[|p=��!cz0|�i�L�;����-�ٕnǺ�-�B%/�=Ŝ�&Q��m��g-�jx�nѨ̵��k�#2ؚ7�b�z�lh�4�̴������^��2Y���nc���1���2�c	z�7��5rR�|�Z�؆5�V�G%��5H�ZJ?���/K���q0�JI��xBG������k�}+I/�I�V�+m!�O����-[>�;�DF�ۗw)2�[A\��~���Ҥ��ah��,UJ�lv�����NS�s�g/Dg{N�=da��`��I*!"�e���jy��/3��v������,]֋o�q�I�?�!��˅��2�=	��6,�ٿy<|���"���?���?ڥ����_&l�/��zz0���d�p�OvGu�����^B�Q��G}�Ó�����畤k���W@�&T�J���-���-��|	���l�Y�?r���aaTJX�F����
0�6�66�^�F�p`T��t�'��������Q�3��gF��>G|>׋`�)�AR�9I7�d%O�*g����`�����jnnPY}7��QK��v���'��UͰ(�E�#ʤT�hom3����{�v��'9W�N��/�Lx�9'�Η��c��o��k��xX��t���w1�{;#W	�V�����x�<K[�-OD��*
�8>�l{�V�����Jb+�g$,�xw�f��y�3���g���Vd�>����#�t��u���|']�h�ZlWGZG�u���^�e��<����N?�������q��������W~D����_���AӖ��{��v�k���R������u��SV�s�����(�o��Í�{��#z@~D��������c��{��#У�p��ǍV0>d�����j�*����#�F��Q���QAx�Q!mT�@"�F�0�Qa<Ψ0>Ĩ�bTHA"�F��Q!mT�@5pm�2*���
h�Bڨv�8��0gTbTH	1*���
h�Bڨ�6*D��
(��� �B
ڨ�6*D��Z?jnT�3*�1*��R�F��Q!mT�@"�F��QAx�Q!mT�@"�F���
�C�
)!F��Q!mT�@"�F��Q!eTdTHA"�F�����\���f?��zz���骩�w�Qnu�������Y����l��"fR(�E��r�-��\v?���~�R�,��f
��}#���aW�w#A�w����H��<�}�H0v�֗��R�t���'x�	���p��]c�[�kdvaw��N�Qd���G=��x}) tuG�p�'tuK��j8���+���W=?���~JO//��V؏
��+u�Q��Ԑ$5��KQ�RCT��p`�J	X��g?!Hj�	������0��T���RCV��.5DKQaR��VjH�J	X�!!Hj�	������0�A����RCVjH�`¥��`�!�Kj���%5Ja'�sq������lɉ̖B`��Zi�˖\������	}e�Pzz1xa�(��~T�Ըl�M�p��	X�qْWj\��)5.[��-���eKmR㲥6��g?!Hj\��)5.[��-���eKmR㲥6�q�R��'d/&\j\��)5.[�K�˖ڤ�eKmR㲥6�qْWj\��)5.[��-���eKmR㲥6�q�R�Ըl�+5.[��-uJ�ɖ�O[?�d�����˗%7���<0���A�\��I�?�d�MM��'���m���u�6/tYq��I���oA]?�c��u���J��4���M�n.�֟ۺ��Y��4yG��$�mT���Ǧ��L�?ڥ���xj~���i��j�>~ɥ�e�����Q��e}t�g�u|V��7>��0ޮL����0O{���\��vI㆖涷Sm�M�V���  �� PK-      ! ߤ�lZ                      [Content_Types].xmlPK-      ! ���   N               �  _rels/.relsPK-      ! �d�Q�   1               �  word/_rels/document.xml.relsPK-      ! �y�	  9               �  word/document.xmlPK-      ! �@�$  �               0  word/theme/theme1.xmlPK-      ! +��k�  �	               �  word/settings.xmlPK-      ! �1��  D               d  word/fontTable.xmlPK-      ! �?�b"  N               `  word/webSettings.xmlPK-      ! *zC9~  �               �  docProps/app.xmlPK-      ! v�>r  �               h   docProps/core.xmlPK-      ! ��*  Sp               #  word/styles.xmlPK      �  h.    